module DiceGame();

endmodule